library verilog;
use verilog.vl_types.all;
entity Cache_vlg_vec_tst is
end Cache_vlg_vec_tst;
