library verilog;
use verilog.vl_types.all;
entity CacheController_vlg_vec_tst is
end CacheController_vlg_vec_tst;
